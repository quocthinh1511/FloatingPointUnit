module tim_phan_nguyen (
input wire[7:0]mu,
input wire[7:0]dau,
input [22:0]a,
output reg [23:0]b,
output reg [22:0]c
);  
always @(mu or a)    
if( dau <= 8'h2B)
case (mu)
7'd0: begin b[23:0]<={(22'b0),1'b1}; c[22:0]<=a[22:0]; end 
7'd1: begin b[23:0]<={(22'b0),1'b1,a[22]}; c[22:0]<={a[21:0],1'b0}; end 
7'd2: begin b[23:0]<={(21'b0),1'b1,a[22:21]}; c[22:0]<={a[20:0],2'b0}; end 
7'd3: begin b[23:0]<={(20'b0),1'b1,a[22:20]}; c[22:0]<={a[19:0],3'b0}; end 
7'd4: begin b[23:0]<={(19'b0),1'b1,a[22:19]}; c[22:0]<={a[18:0],4'b0}; end 
7'd5: begin b[23:0]<={(18'b0),1'b1,a[22:18]}; c[22:0]<={a[17:0],5'b0}; end 
7'd6: begin b[23:0]<={(17'b0),1'b1,a[22:17]}; c[22:0]<={a[16:0],6'b0}; end 
7'd7: begin b[23:0]<={(16'b0),1'b1,a[22:16]}; c[22:0]<={a[15:0],7'b0}; end 
7'd8: begin b[23:0]<={(15'b0),1'b1,a[22:15]}; c[22:0]<={a[14:0],8'b0}; end 
7'd9: begin b[23:0]<={(14'b0),1'b1,a[22:14]}; c[22:0]<={a[13:0],9'b0}; end 
7'd10: begin b[23:0]<={(13'b0),1'b1,a[22:13]}; c[22:0]<={a[12:0],10'b0}; end 
7'd11: begin b[23:0]<={(12'b0),1'b1,a[22:12]}; c[22:0]<={a[11:0],11'b0}; end 
7'd12: begin b[23:0]<={(11'b0),1'b1,a[22:11]}; c[22:0]<={a[10:0],12'b0}; end 
7'd13: begin b[23:0]<={(10'b0),1'b1,a[22:10]}; c[22:0]<={a[9:0],13'b0}; end 
7'd14: begin b[23:0]<={(9'b0),1'b1,a[22:9]}; c[22:0]<={a[8:0],14'b0}; end 
7'd15: begin b[23:0]<={(8'b0),1'b1,a[22:8]}; c[22:0]<={a[7:0],15'b0}; end 
7'd16: begin b[23:0]<={(7'b0),1'b1,a[22:7]}; c[22:0]<={a[6:0],16'b0}; end
7'd17: begin b[23:0]<={(6'b0),1'b1,a[22:6]}; c[22:0]<={a[5:0],17'b0}; end 
7'd18: begin b[23:0]<={(5'b0),1'b1,a[22:5]}; c[22:0]<={a[4:0],18'b0}; end 
7'd19: begin b[23:0]<={(4'b0),1'b1,a[22:4]}; c[22:0]<={a[3:0],19'b0}; end 
7'd20: begin b[23:0]<={(3'b0),1'b1,a[22:3]}; c[22:0]<={a[2:0],20'b0}; end 
7'd21: begin b[23:0]<={(2'b0),1'b1,a[22:2]}; c[22:0]<={a[1:0],21'b0}; end 
7'd22: begin b[23:0]<={(1'b0),1'b1,a[22:1]}; c[22:0]<={a[0],22'b0}; end
7'd23: begin b[23:0]<={1'b1,a[22:0]}; c[22:0]<={23'b0}; end 
default begin b[23:0]<={24'b1}; c[22:0]<={23'b0}; end 
endcase 
else  case (mu)
7'd1: begin b[23:0]<={(24'b0)}; c[22:0]<={1'b1,a[22:1]}; end 
7'd2: begin b[23:0]<={(24'b0)}; c[22:0]<={1'b0,1'b1,a[22:2]}; end 
7'd3: begin b[23:0]<={(24'b0)}; c[22:0]<={2'b0,1'b1,a[22:3]}; end 
7'd4: begin b[23:0]<={(24'b0)}; c[22:0]<={3'b0,1'b1,a[22:4]}; end 
7'd5: begin b[23:0]<={(24'b0)}; c[22:0]<={4'b0,1'b1,a[22:5]}; end 
7'd6: begin b[23:0]<={(24'b0)}; c[22:0]<={5'b0,1'b1,a[22:6]}; end 
7'd7: begin b[23:0]<={(24'b0)}; c[22:0]<={6'b0,1'b1,a[22:7]}; end 
7'd8: begin b[23:0]<={(24'b0)}; c[22:0]<={7'b0,1'b1,a[22:8]}; end 
7'd9: begin b[23:0]<={(24'b0)}; c[22:0]<={8'b0,1'b1,a[22:9]}; end 
7'd10: begin b[23:0]<={(24'b0)}; c[22:0]<={9'b0,1'b1,a[22:10]}; end 
7'd11: begin b[23:0]<={(24'b0)}; c[22:0]<={10'b0,1'b1,a[22:11]}; end 
7'd12: begin b[23:0]<={(24'b0)}; c[22:0]<={11'b0,1'b1,a[22:12]}; end 
7'd13: begin b[23:0]<={(24'b0)}; c[22:0]<={12'b0,1'b1,a[22:13]}; end 
7'd14: begin b[23:0]<={(24'b0)}; c[22:0]<={13'b0,1'b1,a[22:14]}; end 
7'd15: begin b[23:0]<={(24'b0)}; c[22:0]<={14'b0,1'b1,a[22:15]}; end 
7'd16: begin b[23:0]<={(24'b0)}; c[22:0]<={15'b0,1'b1,a[22:16]}; end
7'd17: begin b[23:0]<={(24'b0)}; c[22:0]<={16'b0,1'b1,a[22:17]}; end 
7'd18: begin b[23:0]<={(24'b0)}; c[22:0]<={17'b0,1'b1,a[22:18]}; end 
7'd19: begin b[23:0]<={(24'b0)}; c[22:0]<={18'b0,1'b1,a[22:19]}; end 
7'd20: begin b[23:0]<={(24'b0)}; c[22:0]<={19'b0,1'b1,a[22:20]}; end 
7'd21: begin b[23:0]<={(24'b0)}; c[22:0]<={20'b0,1'b1,a[22:21]}; end 
7'd22: begin b[23:0]<={(24'b0)}; c[22:0]<={21'b0,1'b1,a[22]}; end
7'd23: begin b[23:0]<={24'b0}; c[22:0]<={22'b0,1'b1}; end 
default begin b[23:0]<={24'b0}; c[22:0]<={23'b0}; end 


endcase 
endmodule
module t_tim_phan_nguyen;
	reg [7:0]mu;reg [7:0]dau;
	reg [22:0]a;
        wire [23:0]b;
         wire [22:0]c;
parameter time_out = 100;
	tim_phan_nguyen z(.mu(mu),.dau(dau),.a(a),.b(b),.c(c));
      
initial $monitor($time," so mu %d , %b  , %b ,  %b  ", mu,a,b,c );
	initial begin

	#0 dau=8'h2B; mu=8'b0000_0100; a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_0110;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2B;mu=8'b0000_0111;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1000;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1001;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1010;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1011;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1100;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1101;a=23'b100_0001_1111_0000_0000_0000;
        #10 dau=8'h2D;mu=8'b0000_1110;a=23'b100_0001_1111_0000_0000_0000;
	#10 dau=8'h2D;mu=8'b0000_1111;a=23'b100_0001_1111_0000_0000_0000;
end 
endmodule